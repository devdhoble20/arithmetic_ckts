`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.01.2025 14:54:13
// Design Name: 
// Module Name: dadda16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module dadda16(
    input [15:0] a,
    input [15:0] b,
    output [31:0] m);
    wire [23:0] w1;
    wire [87:0] w2;
    wire [107:0] w3;
    wire [91:0] w4;
    wire [51:0] w5;
    
    wire [32:0] m1;
    // Stage 1 : d = 13
    HA HA1 (b[0]&a[13], b[1]&a[12], w1[0], w1[1]);
    
    FA FA1 (b[0]&a[14], b[1]&a[13], b[2]&a[12], w1[2], w1[3]);
    HA HA2 (b[3]&a[11], b[4]&a[10], w1[4], w1[5]);
    
    FA FA2 (b[0]&a[15], b[1]&a[14], b[2]&a[13], w1[6], w1[7]);
    FA FA3 (b[3]&a[12], b[4]&a[11], b[5]&a[10], w1[8], w1[9]);
    HA HA3 (b[6]&a[9], b[7]&a[8], w1[10], w1[11]);
    
    FA FA4 (b[1]&a[15], b[2]&a[14], b[3]&a[13], w1[12], w1[13]);
    FA FA5 (b[4]&a[12], b[5]&a[11], b[6]&a[10], w1[14], w1[15]);
    HA HA4 (b[7]&a[9], b[8]&a[8], w1[16], w1[17]);
    
    FA FA6 (b[2]&a[15], b[3]&a[14], b[4]&a[13], w1[18], w1[19]);
    FA FA7 (b[5]&a[12], b[6]&a[11], b[7]&a[10], w1[20], w1[21]);
    
    FA FA8 (b[3]&a[15], b[4]&a[14], b[5]&a[13], w1[22], w1[23]);
    
    // Stage 2 : d = 9
    HA HA5 (b[0]&a[9], b[1]&a[8], w2[0], w2[1]);
    
    FA FA9 (b[0]&a[10], b[1]&a[9], b[2]&a[8], w2[2], w2[3]);
    HA HA6 (b[3]&a[7], b[4]&a[6], w2[4], w2[5]);
    
    FA FA10 (b[0]&a[11], b[1]&a[10], b[2]&a[9], w2[6], w2[7]);
    FA FA11 (b[3]&a[8], b[4]&a[7], b[5]&a[6], w2[8], w2[9]);
    HA HA7 (b[6]&a[5], b[7]&a[4], w2[10], w2[11]);
    
    FA FA12 (b[0]&a[12], b[1]&a[11], b[2]&a[10], w2[12], w2[13]);
    FA FA13 (b[3]&a[9], b[4]&a[8], b[5]&a[7], w2[14], w2[15]);
    FA FA14 (b[6]&a[6], b[7]&a[5], b[8]&a[4], w2[16], w2[17]);
    HA HA8 (b[9]&a[3], b[10]&a[2], w2[18], w2[19]);
    
    FA FA15 (w1[0], b[2]&a[11], b[3]&a[10], w2[20], w2[21]);
    FA FA16 (b[4]&a[9], b[5]&a[8], b[6]&a[7], w2[22], w2[23]);
    FA FA17 (b[7]&a[6], b[8]&a[5], b[9]&a[4], w2[24], w2[25]);
    FA FA18 (b[10]&a[3], b[11]&a[2], b[12]&a[1], w2[26], w2[27]);
    
    FA FA19 (w1[2],w1[1],w1[4],w2[28], w2[29]);
    FA FA20 (b[5]&a[9], b[6]&a[8], b[7]&a[7], w2[30], w2[31]);
    FA FA21 (b[8]&a[6], b[9]&a[5], b[10]&a[4], w2[32], w2[33]);
    FA FA22 (b[11]&a[3], b[12]&a[2], b[13]&a[1], w2[34], w2[35]);
    
    FA FA23 (w1[6], w1[3], w1[8], w2[36], w2[37]);
    FA FA24 (w1[10], w1[5], b[8]&a[7], w2[38], w2[39]);
    FA FA25 (b[9]&a[6], b[10]&a[5], b[11]&a[4], w2[40], w2[41]);
    FA FA26 (b[12]&a[3], b[13]&a[2], b[14]&a[1], w2[42], w2[43]);
    
    FA FA27 (w1[12], w1[7], w1[14], w2[44], w2[45]);
    FA FA28 (w1[9], w1[16], w1[11], w2[46], w2[47]);
    FA FA29 (b[9]&a[7], b[10]&a[6], b[11]&a[5], w2[48], w2[49]);
    FA FA30 (b[12]&a[4], b[13]&a[3], b[14]&a[2], w2[50], w2[51]);
    
    FA FA31 (w1[18], w1[13], w1[20], w2[52], w2[53]);
    FA FA32 (w1[15], b[8]&a[9], w1[17], w2[54], w2[55]);
    FA FA33 (b[9]&a[8], b[10]&a[7], b[11]&a[6], w2[56], w2[57]);
    FA FA34 (b[12]&a[5], b[13]&a[4], b[14]&a[3], w2[58], w2[59]);
    
    FA FA35 (w1[22], w1[19], b[6]&a[12], w2[60], w2[61]);
    FA FA36 (w1[21], b[7]&a[11], b[8]&a[10], w2[62], w2[63]);
    FA FA37 (b[9]&a[9], b[10]&a[8], b[11]&a[7], w2[64], w2[65]);
    FA FA38 (b[12]&a[6], b[13]&a[5], b[14]&a[4], w2[66], w2[67]);
    
    FA FA39 (b[4]&a[15], w1[23], b[5]&a[14], w2[68], w2[69]);
    FA FA40 (b[6]&a[13], b[7]&a[12], b[8]&a[11], w2[70], w2[71]);
    FA FA41 (b[9]&a[10], b[10]&a[9], b[11]&a[8], w2[72], w2[73]);
    FA FA42 (b[12]&a[7], b[13]&a[6], b[14]&a[5], w2[74], w2[75]);
    
    FA FA43 (b[5]&a[15], b[6]&a[14], b[7]&a[13], w2[76], w2[77]);
    FA FA44 (b[8]&a[12], b[9]&a[11], b[10]&a[10], w2[78], w2[79]);
    FA FA45 (b[11]&a[9], b[12]&a[8], b[13]&a[7], w2[80], w2[81]);
    
    FA FA46 (b[6]&a[15], b[7]&a[14], b[8]&a[13], w2[82], w2[83]);
    FA FA47 (b[9]&a[12], b[10]&a[11], b[11]&a[10], w2[84], w2[85]);
    
    FA FA48 (b[7]&a[15], b[8]&a[14], b[9]&a[13], w2[86], w2[87]);
    
    // Stage 3 : d = 6
    HA HA9 (b[0]&a[6], b[1]&a[5], w3[0], w3[1]);
    
    FA FA49 (b[0]&a[7], b[1]&a[6], b[2]&a[5], w3[2], w3[3]);
    HA HA10 (b[3]&a[4], b[4]&a[3], w3[4], w3[5]);
    
    FA FA50 (b[0]&a[8], b[1]&a[7], b[2]&a[6], w3[6], w3[7]);
    FA FA51 (b[3]&a[5], b[4]&a[4], b[5]&a[3], w3[8], w3[9]);
    HA HA11 (b[6]&a[2], b[7]&a[1], w3[10], w3[11]);
    
    FA FA52 (w2[0], b[2]&a[7], b[3]&a[6], w3[12], w3[13]);
    FA FA53 (b[4]&a[5], b[5]&a[4], b[6]&a[3], w3[14], w3[15]);
    FA FA54 (b[7]&a[2], b[8]&a[1], b[9]&a[0], w3[16], w3[17]);
    
    FA FA55 (w2[2], w2[1], w2[4], w3[18], w3[19]);
    FA FA56 (b[5]&a[5], b[6]&a[4], b[7]&a[3], w3[20], w3[21]);
    FA FA57 (b[8]&a[2], b[9]&a[1], b[10]&a[0], w3[22], w3[23]);
    
    FA FA58 (w2[6], w2[3], w2[8], w3[24], w3[25]);
    FA FA59 (w2[5], w2[10], b[8]&a[3], w3[26], w3[27]);
    FA FA60 (b[9]&a[2], b[10]&a[1], b[11]&a[0], w3[28], w3[29]);
    
    FA FA61 (w2[12], w2[7], w2[14], w3[30], w3[31]);
    FA FA62 (w2[9], w2[16], w2[11], w3[32], w3[33]);
    FA FA63 (w2[18], b[11]&a[1], b[12]&a[0], w3[34], w3[35]);
    
    FA FA64 (w2[20], w2[13], w2[22], w3[36], w3[37]);
    FA FA65 (w2[24], w2[15], w2[17], w3[38], w3[39]);
    FA FA66 (w2[26], w2[19], b[13]&a[0], w3[40], w3[41]);
    
    FA FA67 (w2[28], w2[30], w2[21], w3[42], w3[43]);
    FA FA68 (w2[32], w2[23], w2[25], w3[44], w3[45]);
    FA FA69 (w2[34], w2[27], b[14]&a[0], w3[46], w3[47]);
    
    FA FA70 (w2[36], w2[29], w2[38], w3[48], w3[49]);
    FA FA71 (w2[31], w2[40], w2[33], w3[50], w3[51]);
    FA FA72 (w2[42], w2[35], b[15]&a[0], w3[52], w3[53]);
    
    FA FA73 (w2[44], w2[37], w2[46], w3[54], w3[55]);
    FA FA74 (w2[48], w2[39], w2[41], w3[56], w3[57]);
    FA FA75 (w2[50], w2[43], b[15]&a[1], w3[58], w3[59]);
    
    FA FA76 (w2[52], w2[45], w2[54], w3[60], w3[61]);
    FA FA77 (w2[47], w2[56], w2[49], w3[62], w3[63]);
    FA FA78 (w2[58], w2[51], b[15]&a[2], w3[64], w3[65]);
    
    FA FA79 (w2[60], w2[53], w2[62], w3[66], w3[67]);
    FA FA80 (w2[55], w2[64], w2[57], w3[68], w3[69]);
    FA FA81 (w2[66], w2[59], b[15]&a[3], w3[70], w3[71]);
    
    FA FA82 (w2[68], w2[61], w2[70], w3[72], w3[73]);
    FA FA83 (w2[63], w2[72], w2[65], w3[74], w3[75]);
    FA FA84 (w2[74], w2[67], b[15]&a[4], w3[76], w3[77]);
    
    FA FA85 (w2[76], w2[69], w2[78], w3[78], w3[79]);
    FA FA86 (w2[71], w2[80], w2[73], w3[80], w3[81]);
    FA FA87 (b[14]&a[6], w2[75], b[15]&a[5], w3[82], w3[83]);
    
    FA FA88 (w2[82], w2[77], w2[84], w3[84], w3[85]);
    FA FA89 (w2[79], w2[81], b[12]&a[9], w3[86], w3[87]);
    FA FA90 (b[13]&a[8], b[14]&a[7], b[15]&a[6], w3[88], w3[89]);
    
    FA FA91 (w2[86], w2[83], b[10]&a[12], w3[90], w3[91]);
    FA FA92 (w2[85], b[11]&a[11], b[12]&a[10], w3[92], w3[93]);
    FA FA93 (b[13]&a[9], b[14]&a[8], b[15]&a[7], w3[94], w3[95]);
    
    FA FA94 (b[8]&a[15], w2[87], b[9]&a[14], w3[96], w3[97]);
    FA FA95 (b[10]&a[13], b[11]&a[12], b[12]&a[11], w3[98], w3[99]);
    FA FA96 (b[13]&a[10], b[14]&a[9], b[15]&a[8], w3[100], w3[101]);
    
    FA FA97 (b[9]&a[15], b[10]&a[14], b[11]&a[13], w3[102], w3[103]);
    FA FA98 (b[12]&a[12], b[13]&a[11], b[14]&a[10], w3[104], w3[105]);
    
    FA FA99 (b[10]&a[15], b[11]&a[14], b[12]&a[13], w3[106], w3[107]);
    
    // Stage 4 : d = 4
    HA HA12 (b[0]&a[4], b[1]&a[3], w4[0], w4[1]);
    
    FA FA100 (b[0]&a[5], b[1]&a[4], b[2]&a[3], w4[2], w4[3]);
    HA HA13 (b[3]&a[2], b[4]&a[1], w4[4], w4[5]);
    
    FA FA101 (w3[0], b[2]&a[4], b[3]&a[3], w4[6], w4[7]);
    FA FA102 (b[4]&a[2], b[5]&a[1], b[6]&a[0], w4[8], w4[9]);
    
    FA FA103 (w3[2], w3[1], w3[4], w4[10], w4[11]);
    FA FA104 (b[5]&a[2], b[6]&a[1], b[7]&a[0], w4[12], w4[13]);
    
    FA FA105 (w3[6], w3[8], w3[3], w4[14], w4[15]);
    FA FA106 (w3[5], w3[10], b[8]&a[0], w4[16], w4[17]);
    
    FA FA107 (w3[12], w3[14], w3[7], w4[18], w4[19]);
    FA FA108 (w3[9], w3[16], w3[11], w4[20], w4[21]);
    
    FA FA109 (w3[18], w3[13], w3[20], w4[22], w4[23]);
    FA FA110 (w3[15], w3[22], w3[17], w4[24], w4[25]);
    
    FA FA111 (w3[24], w3[26], w3[19], w4[26], w4[27]);
    FA FA112 (w3[21], w3[28], w3[23], w4[28], w4[29]);
    
    FA FA113 (w3[30], w3[25], w3[32], w4[30], w4[31]);
    FA FA114 (w3[27], w3[34], w3[29], w4[32], w4[33]);
    
    FA FA115 (w3[36], w3[38], w3[31], w4[34], w4[35]);
    FA FA116 (w3[33], w3[40], w3[35], w4[36], w4[37]);
    
    FA FA117 (w3[42], w3[37], w3[44], w4[38], w4[39]);
    FA FA118 (w3[39], w3[46], w3[41], w4[40], w4[41]);
    
    FA FA119 (w3[48], w3[43], w3[50], w4[42], w4[43]);
    FA FA120 (w3[45], w3[52], w3[47], w4[44], w4[45]);
    
    FA FA121 (w3[54], w3[49], w3[56], w4[46], w4[47]);
    FA FA122 (w3[51], w3[58], w3[53], w4[48], w4[49]);
    
    FA FA123 (w3[60], w3[62], w3[55], w4[50], w4[51]);
    FA FA124 (w3[57], w3[64], w3[59], w4[52], w4[53]);
    
    FA FA125 (w3[66], w3[61], w3[68], w4[54], w4[55]);
    FA FA126 (w3[63], w3[70], w3[65], w4[56], w4[57]);
    
    FA FA127 (w3[72], w3[67], w3[74], w4[58], w4[59]);
    FA FA128 (w3[69], w3[76], w3[71], w4[60], w4[61]);
    
    FA FA129 (w3[78], w3[80], w3[73], w4[62], w4[63]);
    FA FA130 (w3[75], w3[82], w3[77], w4[64], w4[65]);
    
    FA FA131 (w3[84], w3[79], w3[86], w4[66], w4[67]);
    FA FA132 (w3[81], w3[88], w3[83], w4[68], w4[69]);
    
    FA FA133 (w3[90], w3[85], w3[92], w4[70], w4[71]);
    FA FA134 (w3[87], w3[94], w3[89], w4[72], w4[73]);
    
    FA FA135 (w3[96], w3[91], w3[98], w4[74], w4[75]);
    FA FA136 (w3[93], w3[100], w3[95], w4[76], w4[77]);
    
    FA FA137 (w3[102], w3[97], w3[104], w4[78], w4[79]);
    FA FA138 (w3[101], b[15]&a[9], w3[99], w4[80], w4[81]);
    
    FA FA139 (w3[106], w3[103], b[13]&a[12], w4[82], w4[83]);
    FA FA140 (b[14]&a[11], b[15]&a[10], w3[105], w4[84], w4[85]);
    
    FA FA141 (b[11]&a[15], w3[107], b[12]&a[14], w4[86], w4[87]);
    FA FA142 (b[13]&a[13], b[14]&a[12], b[15]&a[11], w4[88], w4[89]);
    
    FA FA143 (b[12]&a[15], b[13]&a[14], b[14]&a[13], w4[90], w4[91]);
    
    // Stage 5 : d = 3
    HA HA14 (b[0]&a[3], b[1]&a[2], w5[0], w5[1]);
    
    FA FA144 (w4[0], b[2]&a[2], b[3]&a[1], w5[2], w5[3]);
    
    FA FA145 (w4[2], w4[1], w4[4], w5[4], w5[5]);
    
    FA FA146 (w4[6], w4[3], w4[8], w5[6], w5[7]);
    
    FA FA147 (w4[10], w4[7], w4[12], w5[8], w5[9]);
    
    FA FA148 (w4[14], w4[11], w4[16], w5[10], w5[11]);
    
    FA FA149 (w4[18], w4[15], w4[20], w5[12], w5[13]);
    
    FA FA150 (w4[22], w4[19], w4[24], w5[14], w5[15]);
    
    FA FA151 (w4[26], w4[23], w4[28], w5[16], w5[17]);
    
    FA FA152 (w4[30], w4[27], w4[32], w5[18], w5[19]);
    
    FA FA153 (w4[34], w4[31], w4[36], w5[20], w5[21]);
    
    FA FA154 (w4[38], w4[35], w4[40], w5[22], w5[23]);
    
    FA FA155 (w4[42], w4[39], w4[44], w5[24], w5[25]);
    
    FA FA156 (w4[46], w4[43], w4[48], w5[26], w5[27]);
    
    FA FA157 (w4[50], w4[47], w4[52], w5[28], w5[29]);
    
    FA FA158 (w4[54], w4[51], w4[56], w5[30], w5[31]);
    
    FA FA159 (w4[58], w4[55], w4[60], w5[32], w5[33]);
    
    FA FA160 (w4[62], w4[59], w4[64], w5[34], w5[35]);
    
    FA FA161 (w4[66], w4[63], w4[68], w5[36], w5[37]);
    
    FA FA162 (w4[70], w4[67], w4[72], w5[38], w5[39]);
    
    FA FA163 (w4[74], w4[71], w4[76], w5[40], w5[41]);
    
    FA FA164 (w4[78], w4[75], w4[80], w5[42], w5[43]);
    
    FA FA165 (w4[82], w4[79], w4[84], w5[44], w5[45]);
    
    FA FA166 (w4[86], w4[83], w4[88], w5[46], w5[47]);
    
    FA FA167 (w4[90], w4[87], b[15]&a[12], w5[48], w5[49]);
    
    FA FA168 (b[13]&a[15], w4[91], b[14]&a[14], w5[50], w5[51]);
    
    // Stage 6 : d = 2
    wire [27:0] w6;
    wire [27:0] w7;
    
    HA HA15 (b[0]&a[2], b[1]&a[1], w6[0], w7[0]);
    
    FA FA169 (w5[0], b[2]&a[1], b[3]&a[0], w6[1], w7[1]);
    
    FA FA170 (w5[2], w5[1], b[4]&a[0], w6[2], w7[2]);
    
    FA FA171 (w5[4], w5[3], b[5]&a[0], w6[3], w7[3]);
    
    FA FA172 (w5[6], w5[5], w4[5], w6[4], w7[4]);
    
    FA FA173 (w5[8], w5[7], w4[9], w6[5], w7[5]);
    
    FA FA174 (w5[10], w5[9], w4[13], w6[6], w7[6]);
    
    FA FA175 (w5[12], w5[11], w4[17], w6[7], w7[7]);
    
    FA FA176 (w5[14], w5[13], w4[21], w6[8], w7[8]);
    
    FA FA177 (w5[16], w5[15], w4[25], w6[9], w7[9]);
    
    FA FA178 (w5[18], w5[17], w4[29], w6[10], w7[10]);
    
    FA FA179 (w5[20], w5[19], w4[33], w6[11], w7[11]);
    
    FA FA180 (w5[22], w5[21], w4[37], w6[12], w7[12]);
    
    FA FA181 (w5[24], w5[23], w4[41], w6[13], w7[13]);
    
    FA FA182 (w5[26], w5[25], w4[45], w6[14], w7[14]);
    
    FA FA183 (w5[28], w5[27], w4[49], w6[15], w7[15]);
    
    FA FA184 (w5[30], w5[29], w4[53], w6[16], w7[16]);
    
    FA FA185 (w5[32], w5[31], w4[57], w6[17], w7[17]);
    
    FA FA186 (w5[34], w5[33], w4[61], w6[18], w7[18]);
    
    FA FA187 (w5[36], w5[35], w4[65], w6[19], w7[19]);
    
    FA FA188 (w5[38], w5[37], w4[69], w6[20], w7[20]);
    
    FA FA189 (w5[40], w5[39], w4[73], w6[21], w7[21]);
    
    FA FA190 (w5[42], w5[41], w4[77], w6[22], w7[22]);
    
    FA FA191 (w5[44], w5[43], w4[81], w6[23], w7[23]);
    
    FA FA192 (w5[46], w5[45], w4[85], w6[24], w7[24]);
    
    FA FA193 (w5[48], w5[47], w4[89], w6[25], w7[25]);
    
    FA FA194 (w5[50], w5[49], b[15]&a[13], w6[26], w7[26]);
    
    FA FA195 (b[14]&a[15], b[15]&a[14], w5[51], w6[27], w7[27]);
    
    // Fast Adder (BK Adder) 
    
    bkadder bk ({0, 0, b[15]&a[15], w6, b[0]&a[1]}, {0, 0, w7, b[2]&a[0], b[1]&a[0]}, 0, m1[31:0], m1[32]);
    assign m[0] = a[0]&b[0];
    assign m[31:1] = m1[30:0];
    
endmodule

module HA(input x, input y, output s, output c);
    assign s = x^y;
    assign c = x&y;
endmodule

module FA(input x, input y, input z, output s, output c);
    assign s = x^y^z;
    assign c = (x&y) | (y&z) | (z&x);
endmodule
